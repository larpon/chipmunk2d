// Copyright(C) 2025 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module chipmunk2d

//
// cpTransform.h
//

// TODO Non-numerical: #define CHIPMUNK_TRANSFORM_H
